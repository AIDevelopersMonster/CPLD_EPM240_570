// ============================================================
// Имя файла: my_uart_rx.v
// Описание: Модуль для приема данных по UART (RS232).
//           Обрабатывает входящие данные, синхронизирует их по скорости передачи данных,
//           генерирует сигнал прерывания при получении данных и готовит данные для дальнейшей обработки.
//           Модуль генерирует тактовые сигналы для приема данных и синхронизирует их с тактовым сигналом.
//
// Создано: AIDevelopersMonster
// Репозиторий GitHub: https://github.com/AIDevelopersMonster/CPLD_EPM240_570/
//
// ============================================================


`timescale 1ns / 1ps

module my_uart_rx(
				clk,rst_n,
				rs232_rx,rx_data,rx_int,
				clk_bps,bps_start
			);

input clk;		// Входной тактовый сигнал 50MHz
input rst_n;	// Низкий активный сигнал сброса
input rs232_rx;	// Входной сигнал для приема данных по RS232
input clk_bps;	// Тактовый сигнал для синхронизации передачи данных (baud rate)
output bps_start;		// Сигнал начала передачи для синхронизации
output[7:0] rx_data;	// Принятые 8 бит данных
output rx_int;	// Сигнал прерывания для уведомления о начале приема данных

//----------------------------------------------------------------
// Регистры для сдвига входных данных
//----------------------------------------------------------------
reg rs232_rx0, rs232_rx1, rs232_rx2, rs232_rx3;  // Сдвиговые регистры для приема
wire neg_rs232_rx;  // Сигнал для обнаружения переднего фронта

// Процесс сдвига данных для корректной синхронизации
always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        rs232_rx0 <= 1'b0;
        rs232_rx1 <= 1'b0;
        rs232_rx2 <= 1'b0;
        rs232_rx3 <= 1'b0;
    end else begin
        rs232_rx0 <= rs232_rx;
        rs232_rx1 <= rs232_rx0;
        rs232_rx2 <= rs232_rx1;
        rs232_rx3 <= rs232_rx2;
    end
end

// Обнаружение переднего фронта сигнала приема (RS232)
assign neg_rs232_rx = rs232_rx3 & rs232_rx2 & ~rs232_rx1 & ~rs232_rx0;  // Сигнал для старта приема

//----------------------------------------------------------
// Логика для управления сигналом начала передачи и прерывания
//----------------------------------------------------------

reg bps_start_r;
reg [3:0] num;  // Счетчик для отслеживания приема битов данных
reg rx_int;      // Сигнал прерывания для уведомления о получении данных

// Процесс для генерации сигнала начала передачи и прерывания
always @ (posedge clk or negedge rst_n)
    if (!rst_n) begin
        bps_start_r <= 1'bz;
        rx_int <= 1'b0;
    end else if (neg_rs232_rx) begin  // Если был обнаружен передний фронт сигнала
        bps_start_r <= 1'b1;           // Начало передачи данных
        rx_int <= 1'b1;                // Генерация прерывания для приема данных
    end else if (num == 4'd11) begin  // Если 11 бит принято (старт + 8 данных + стоп)
        bps_start_r <= 1'b0;           // Завершение передачи
        rx_int <= 1'b0;                // Отключение прерывания
    end

assign bps_start = bps_start_r;  // Выходной сигнал начала передачи

//----------------------------------------------------------
// Регистры для хранения данных
//----------------------------------------------------------

reg [7:0] rx_data_r;  // Принятый байт данных
reg [7:0] rx_temp_data;  // Временный регистр для данных

// Процесс приема данных по битам
always @ (posedge clk or negedge rst_n)
    if (!rst_n) begin
        rx_temp_data <= 8'd0;
        num <= 4'd0;
        rx_data_r <= 8'd0;
    end else if (rx_int) begin  // Если активен сигнал прерывания
        if (clk_bps) begin  // Прием данных по тактовому сигналу
            num <= num + 1'b1;
            case (num)
                4'd1: rx_temp_data[0] <= rs232_rx;  // Прием бита 0
                4'd2: rx_temp_data[1] <= rs232_rx;  // Прием бита 1
                4'd3: rx_temp_data[2] <= rs232_rx;  // Прием бита 2
                4'd4: rx_temp_data[3] <= rs232_rx;  // Прием бита 3
                4'd5: rx_temp_data[4] <= rs232_rx;  // Прием бита 4
                4'd6: rx_temp_data[5] <= rs232_rx;  // Прием бита 5
                4'd7: rx_temp_data[6] <= rs232_rx;  // Прием бита 6
                4'd8: rx_temp_data[7] <= rs232_rx;  // Прием бита 7
                default: ;
            endcase
        end else if (num == 4'd11) begin  // Если все 11 бит принято (старт + 8 данных + стоп)
            num <= 4'd0;                     // Сброс счетчика
            rx_data_r <= rx_temp_data;       // Перенос данных в основной регистр
        end
    end

assign rx_data = rx_data_r;  // Выходной сигнал с принятыми данными

endmodule