/*
  --------------------------------------------------------------------------------
  Модуль     : led_twinkle.v
  Описание   : Этот модуль генерирует эффект мигания для 8-битного вывода LED.
                Светодиод переключается каждую секунду в зависимости от входного
                тактового сигнала 50 МГц.
  
  Автор      : kontakts.ru
  Дата       : 21-10-2023
  
  Файл       : led_twinkle.v
  Язык       : Verilog
  
  Лицензия   : Open-source (указать лицензию, если необходимо)
  --------------------------------------------------------------------------------
*/

/*
  Модуль использует входной тактовый сигнал 50 МГц (`clk`) и генерирует 8-битный
  выход (`led`). Состояние светодиода переключается каждые 25 миллионов тактовых
  циклов, что соответствует примерно одной секунде (при тактовой частоте 50 МГц).
  
  Счётчик увеличивается на каждом такте, и когда он достигает значения в 25 миллионов,
  состояние светодиода переключается, а счётчик сбрасывается.
*/

module led_twinkle(led, clk);  // Определение модуля: "led_twinkle" управляет 8-битным светодиодом
  
  // Входные и выходные сигналы
  input clk;                  // Входной тактовый сигнал (50 МГц)
  output [8:1] led;           // 8-битный выход для управления светодиодом (1 байт)
  
  // Внутренние регистры
  reg [8:1] led;              // Регистр для хранения состояния светодиода (8 бит)
  reg [24:0] counter;         // 25-битный счётчик для отслеживания тактовых циклов
  
  /*
    Блок Always: Срабатывает при каждом положительном фронте тактового сигнала.
    Этот блок отслеживает количество тактов и переключает светодиод, когда счётчик
    достигает значения, соответствующего 1 секунде (25 миллионов тактов).
  */
  always @(posedge clk) begin
    counter <= counter + 1;  // Увеличиваем счётчик на каждом тактовом цикле
    
    // Когда счётчик достигает 25 миллионов (1 секунда), переключаем светодиод и сбрасываем счётчик
    if (counter == 25'd25000000) begin
      led <= ~led;           // Переключаем состояние светодиода (инвертируем биты)
      counter <= 0;          // Сбрасываем счётчик после переключения светодиода
    end
  end
  
endmodule
