/*******************************************************************
** FPGA проект - Скрипт для управления семисегментным дисплеем
** Вебсайт: www.kontakts.ru
** Магазин: 
** Контакт: 
** Этот код предназначен для использования с FPGA для динамического
** отображения чисел на семисегментном дисплее, используя алгоритм сканирования.
** Версия: 1.1
** Дата: 01.06.2026
**
** Описание:
** Этот модуль управляет семисегментным дисплеем, сканируя 8 разрядов и отображая
** на них 32-битные данные. Модуль использует 1кГц тактовый сигнал для обновления
** дисплея. Каждое число на дисплее отображается поочередно в течение каждого такта.
** Для изменения частоты можно подстроить значения F_DIV и F_DIV_WIDTH.
*********************************************************************/

module scan_led(clk_1k, d, dig, seg);  // Модуль scan_led для управления семисегментным дисплеем

input clk_1k;          // Входной тактовый сигнал 1 кГц
input [31:0] d;        // Данные, которые нужно отобразить (32 бита)
output [7:0] dig;      // Выход, определяющий, какой из 8 разрядов активен
output [7:0] seg;      // Выход для семисегментного дисплея

// Регистры для хранения состояний сегментов и разрядов
reg [7:0] seg_r;       // Регистр для отображения сегментов
reg [7:0] dig_r;       // Регистр для выбора активного разряда
reg [3:0] disp_dat;    // Регистр для хранения данных для отображения
reg [2:0] count;       // Счётчик для выборки разрядов

// Присваивание выходных значений
assign dig = dig_r;    // Назначение состояния разрядов
assign seg = seg_r;    // Назначение состояния сегментов

// Счётчик для обновления дисплея каждый такт
always @(posedge clk_1k) 
begin
    count <= count + 1'b1;  // Увеличиваем счётчик на каждом такте
end

// Выбор данных для отображения в зависимости от состояния счётчика
always @(posedge clk_1k) 
begin
    case(count)   // Выбор разряда для отображения
        3'd0: disp_dat = d[31:28];  // Отображение первых 4 бит
        3'd1: disp_dat = d[27:24];  // Отображение следующих 4 бит
        3'd2: disp_dat = d[23:20];  // И так далее
        3'd3: disp_dat = d[19:16];
        3'd4: disp_dat = d[15:12];
        3'd5: disp_dat = d[11:8];
        3'd6: disp_dat = d[7:4];
        3'd7: disp_dat = d[3:0];
    endcase
    
    // Настройка активации разряда
    case(count)
        3'd0: dig_r = 8'b01111111;  // Активация первого разряда
        3'd1: dig_r = 8'b10111111;  // Активация второго разряда
        3'd2: dig_r = 8'b11011111;  // Активация третьего разряда
        3'd3: dig_r = 8'b11101111;  // Активация четвёртого разряда
        3'd4: dig_r = 8'b11110111;  // Активация пятого разряда
        3'd5: dig_r = 8'b11111011;  // Активация шестого разряда
        3'd6: dig_r = 8'b11111101;  // Активация седьмого разряда
        3'd7: dig_r = 8'b11111110;  // Активация восьмого разряда
    endcase    
end

// Отображение символов на дисплее в зависимости от данных
always @(disp_dat)
begin
    case(disp_dat)  // Сопоставление данных с сегментами
        4'h0: seg_r = 8'hc0;  // Отображение 0
        4'h1: seg_r = 8'hf9;  // Отображение 1
        4'h2: seg_r = 8'ha4;  // Отображение 2
        4'h3: seg_r = 8'hb0;  // Отображение 3
        4'h4: seg_r = 8'h99;  // Отображение 4
        4'h5: seg_r = 8'h92;  // Отображение 5
        4'h6: seg_r = 8'h82;  // Отображение 6
        4'h7: seg_r = 8'hf8;  // Отображение 7
        4'h8: seg_r = 8'h80;  // Отображение 8
        4'h9: seg_r = 8'h90;  // Отображение 9
        4'ha: seg_r = 8'h88;  // Отображение A
        4'hb: seg_r = 8'h83;  // Отображение B
        4'hc: seg_r = 8'hc6;  // Отображение C
        4'hd: seg_r = 8'ha1;  // Отображение D
        4'he: seg_r = 8'h86;  // Отображение E
        4'hf: seg_r = 8'h8e;  // Отображение F
    endcase
end

endmodule
