/*
  Module     : beep_with_ckey_pins_pnp.v
  Created By : kontakts.ru
  Description: Модуль генерации звукового сигнала с использованием ползунков ckey[1] ~ ckey[4].
               Ползунок ckey[4] управляет включением/выключением зуммера, остальные ползунки включают зуммер с различными эффектами.
               Управление PNP транзистором, база которого подтянута к питанию.
*/

module beep (
    input clk,            // Входной тактовый сигнал (например, 50 МГц)
    input [4:1] ckey,     // Входной сигнал ползунков (ckey[1] ~ ckey[4])
    output beep           // Выходной сигнал для звукового устройства (например, динамик)
);

// Регистр для хранения состояния звукового сигнала
reg beep_r;              // Состояние сигнала
// Регистр для счётчика, который делит частоту входного тактового сигнала
reg [27:0] count;        // Счётчик (длина счётчика зависит от требуемой частоты)

// Логика включения/выключения зуммера
// Инвертируем сигнал для управления PNP транзистором
assign beep = (ckey[4]) ? 1'b1 : ~beep_r; // Если ckey[4] включен, зуммер выключен

// Синхронизация счётчика с тактовым сигналом
always @(posedge clk) begin
    count <= count + 1'b1; // Увеличение счётчика при каждом тактовом импульсе
end

// Логика генерации звукового сигнала
always @(count[9] or ckey[1] or ckey[2] or ckey[3] or ckey[4]) begin
    if (ckey[4] == 1) begin
        beep_r = 1'b0; // Зуммер выключен, если ckey[4] включен
    end else begin
        // Включение зуммера с разными эффектами в зависимости от ckey[1], ckey[2], ckey[3]
        if (ckey[1] == 1) begin
            beep_r = !(count[13] & count[24] & count[27]); // Эффект для ckey[1]
        end else if (ckey[2] == 1) begin 
    beep_r = !(count[15]); // ПРОСТО МЕАНДР 763 Гц
end else if (ckey[3] == 1) begin
    beep_r = !(count[17]); // ПРОСТО МЕАНДР 191 Гц
end else begin
            beep_r = 1'b0; // Если все ползунки выключены, зуммер не работает
        end
    end
end

endmodule