/*******************************************************************
** FPGA проект - Генерация частоты с заданным делителем
** Вебсайт: 
** Магазин: 
** Контакт: 
** Описание:
** Этот модуль генерирует выходной тактовый сигнал с частотой,
** определяемой делителем входного сигнала clock. 
** Частота делителя задается параметром F_DIV, а ширина делителя 
** - параметром F_DIV_WIDTH.
** Процесс деления используется для создания сигнала с 
** 50%-ным скважином и частотой в зависимости от F_DIV.
** Версия: 1.1
** Дата: 01.06.2026
*********************************************************************/

module int_div(clock, clk_out);  // Модуль для делителя частоты

// Входные/выходные сигналы
input clock;        // Входной тактовый сигнал
output clk_out;     // Выходной тактовый сигнал с делённой частотой

// Регистр для хранения состояния сигнала
reg clk_p_r;        // Регистры для положительного и отрицательного сигнала
reg clk_n_r;        
reg [F_DIV_WIDTH - 1:0] count_p;  // Счётчики для деления
reg [F_DIV_WIDTH - 1:0] count_n;

// Параметры делителя
parameter F_DIV = 48000000;  // Частота делителя (можно изменить)
parameter F_DIV_WIDTH = 32;  // Ширина счётчика делителя

// Сигналы флагов деления
wire full_div_p;    // Флаг полного деления для положительного сигнала
wire half_div_p;    // Флаг половинного деления для положительного сигнала
wire full_div_n;    // Флаг полного деления для отрицательного сигнала
wire half_div_n;    // Флаг половинного деления для отрицательного сигнала

// Логика деления (подсчёт делений)
assign full_div_p = (count_p < F_DIV - 1);
assign half_div_p = (count_p < (F_DIV >> 1) - 1);
assign full_div_n = (count_n < F_DIV - 1);
assign half_div_n = (count_n < (F_DIV >> 1) - 1);

// Генерация выходного сигнала
assign clk_out = (F_DIV == 1) ? clock : (F_DIV[0] ? (clk_p_r & clk_n_r) : clk_p_r);

// Логика для положительного делителя
always @(posedge clock) 
begin
    if(full_div_p) 
    begin
        count_p <= count_p + 1'b1;  // Увеличиваем счётчик для положительного сигнала
        if(half_div_p)
            clk_p_r <= 1'b0;   // Если половина делителя, сигнал 0
        else
            clk_p_r <= 1'b1;   // В противном случае, сигнал 1
    end
    else
    begin
        count_p <= 0;   // Сброс счётчика
        clk_p_r <= 1'b0; // Сброс положительного сигнала
    end
end

// Логика для отрицательного делителя
always @(negedge clock) 
begin
    if(full_div_n) 
    begin
        count_n <= count_n + 1'b1;  // Увеличиваем счётчик для отрицательного сигнала
        if(half_div_n)
            clk_n_r <= 1'b0;   // Если половина делителя, сигнал 0
        else
            clk_n_r <= 1'b1;   // В противном случае, сигнал 1
    end
    else
    begin
        count_n <= 0;   // Сброс счётчика
        clk_n_r <= 1'b0; // Сброс отрицательного сигнала
    end
end

endmodule
