// Однострочный комментарий в Verilog начинается с символов // 
// Многострочные комментарии начинаются с /* и заканчиваются на */.

/*
  Модуль    : ckey_led.v
  Автор     : kontakts.ru
  Дата создания : 25-10-2023
*/

module ckey_led( // Имя модуля 'ckey_led' используется для идентификации модуля. 
                // Входные и выходные порты модуля перечисляются ниже.

  input  [MSB_reg:1] ckey,  // Входной сигнал ckey, состоящий из 4 бит (ckey[1] ~ ckey[4])
  output [1:4] led         // Выходной сигнал led, состоящий из 4 бит (led[1] ~ led[4])

);
// Параметр MSB_reg определяет старший разряд для входного сигнала ckey
parameter MSB_reg = 4;

// Присваивание значений между входом и выходом. В данном случае вывод ckey напрямую передается на вывод led.
// В случае с ползунковым переключателем `ckey`, его положение будет напрямую управлять состоянием светодиодов.
// Операция assign используется для назначения значений сигналам и проводникам в Verilog. 
// Эта операция также используется в моделировании потока данных (Data Flow Modeling).
assign led = ckey; 

endmodule

/*
Описание синтаксиса присваивания:
Модуль начинается с ключевого слова module, за которым следует имя модуля и список его входов и выходов. 
Входы и выходы обозначаются с помощью ключевых слов input и output. 

После определения входов и выходов идет описание параметров, переменных и основной логики работы модуля.

В Verilog присваивание значений осуществляется с помощью оператора assign. Этот оператор позволяет передавать значение на сигнал или комбинацию сигналов.
Дополнительно можно использовать параметры "сила передачи" (drive strength) и задержку, но они применяются в основном для моделирования потоков данных, а не для синтеза в реальное оборудование.
*/
