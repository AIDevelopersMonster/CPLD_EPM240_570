// ============================================================
// Имя файла: my_uart_top.v
// Описание: Топ-уровневый модуль для UART-коммуникации.
//           Обрабатывает передачу и прием данных через RS232.
//           Включает обработку данных RX и TX, а также генерацию
//           тактовых сигналов для синхронизации скорости передачи данных (baud rate).
//
// Создано: AIDevelopersMonster
// Репозиторий GitHub: https://github.com/AIDevelopersMonster/CPLD_EPM240_570/
//
// ============================================================

// >>> Директива компилятора: задает единицу времени (1ns) и точность округления (1ps)
// >>> Это важно для симуляции, чтобы понимать реальные временные задержки.
`timescale 1ns / 1ps

module my_uart_top(
    input clk,          // Входной тактовый сигнал 50MHz
    input rst_n,        // Низкий активный сигнал сброса (0 = сброс, 1 = работа)
    input rs232_rx,     // Входной сигнал приема данных RS232 (физический пин)
    output rs232_tx     // Выходной сигнал передачи данных RS232 (физический пин)
);

// ----------------------------------------------------
// Внутренние связи (Wires)
// >>> В Verilog "wire" работает как реальный электрический провод.
// >>> Они не хранят значения, а просто передают сигнал от выхода одного модуля ко входу другого.
// ----------------------------------------------------
wire bps_start1, bps_start2;  // Флаги старта для генераторов частоты (baud rate generators)
wire clk_bps1, clk_bps2;      // Импульсы, указывающие на середину бита данных (для выборки)
wire [7:0] rx_data;           // 8-битная шина данных: передает байт от приемника к передатчику
wire rx_int;                  // Флаг "Прерывание": становится '1', когда приемник закончил получение байта

// ----------------------------------------------------
// Экземпляризация модулей (Instantiation)
// >>> Здесь мы создаем "экземпляры" других модулей и подключаем их к проводам выше.
// ----------------------------------------------------

// 1. Генератор скорости для Приемника (RX)
speed_select speed_rx(
    .clk(clk),           // Системные часы (общие для всех)
    .rst_n(rst_n),       // Общий сброс
    .bps_start(bps_start1), // Вход: сигнал от my_uart_rx, говорящий "начали прием"
    .clk_bps(clk_bps1)      // Выход: тактовый импульс для захвата битов
);

// 2. Модуль Приемника (RX)
my_uart_rx my_uart_rx(
    .clk(clk),
    .rst_n(rst_n),
    .rs232_rx(rs232_rx),    // Вход данных извне
    .rx_data(rx_data),      // Выход: полученный байт данных (идет на вход TX, делая эхо-систему)
    .rx_int(rx_int),        // Выход: сигнал "байт готов" (запускает передачу в TX)
    .clk_bps(clk_bps1),     // Вход: синхроимпульс от speed_select
    .bps_start(bps_start1)  // Выход: управление генератором частоты
);

// 3. Генератор скорости для Передатчика (TX)
speed_select speed_tx(
    .clk(clk),
    .rst_n(rst_n),
    .bps_start(bps_start2), // Вход: сигнал от my_uart_tx
    .clk_bps(clk_bps2)      // Выход: тактовый импульс для отправки битов
);

// 4. Модуль Передатчика (TX)
// >>> Логика работы: Модуль берет данные (rx_data), которые только что пришли,
// >>> и отправляет их обратно (rs232_tx) по сигналу rx_int. Это "Эхо-сервер".
my_uart_tx my_uart_tx(
    .clk(clk),
    .rst_n(rst_n),
    .rx_data(rx_data),      // Вход: данные, полученные от RX
    .rx_int(rx_int),        // Вход: триггер старта передачи (как только RX закончил, TX начинает)
    .rs232_tx(rs232_tx),    // Выход данных наружу
    .clk_bps(clk_bps2),
    .bps_start(bps_start2)
);

endmodule
