//**************************************************************
//  Module     : scan_led.v
//  Created By : (оригинальный автор из китайского примера)
//  Commented  : kontakts.ru
//  Description:
//      Модуль динамической индикации для 8-разрядного 
//      семисегментного индикатора.
//
//      На вход подаётся 32-битное число d, которое интерпретируется
//      как 8 шестнадцатеричных цифр:
//          d[31:28] – старшая цифра (левый разряд),
//          ...
//          d[3:0]   – младшая цифра (правый разряд).
//
//      Модуль поочерёдно включает каждый из 8 разрядов (dig)
//      и выводит соответствующую цифру на сегменты (seg),
//      создавая эффект постоянного свечения за счёт быстрого
//      мультиплексирования.
//
//      clk_1k – тактирование сканирования, обычно ~1 кГц.
//**************************************************************

module scan_led(
    clk_1k,     // тактовый сигнал для сканирования индикатора (~1 кГц)
    d,          // 32-битные данные для отображения (8 hex-цифр)
    dig,        // сигналы выбора разрядов индикатора (аноды/катоды)
    seg         // линии сегментов a..g + точка
);

input        clk_1k;      // входной тактовый сигнал для сканирования
input [31:0] d;           // число, которое нужно вывести (8 * 4 бита)

output [7:0] dig;         // выбор разряда (какой из 8 сейчас активен)
output [7:0] seg;         // шаблон сегментов для выбранного разряда

// Внутренние регистры для выходов
reg [7:0] seg_r;          // текущий шаблон сегментов
reg [7:0] dig_r;          // текущий выбор разряда
reg [3:0] disp_dat;       // 4-битное значение текущей выводимой цифры (0..F)
reg [2:0] count;          // счётчик текущего разряда (0..7)

// Присваиваем регистры внешним выводам
assign dig = dig_r;
assign seg = seg_r;

//--------------------------------------------------------------
// Счётчик разрядов: каждые clk_1k переход по следующему разряду
//--------------------------------------------------------------
always @(posedge clk_1k)
begin
    count <= count + 1'b1;   // 0→1→2→...→7→0→...
end

//--------------------------------------------------------------
// Выбор, какую цифру и какой разряд сейчас отображать
//--------------------------------------------------------------
always @(posedge clk_1k)
begin
    // Выбор 4-битного куска из d в зависимости от count
    case(count)
        3'd0: disp_dat = d[31:28];  // самый левый разряд
        3'd1: disp_dat = d[27:24];
        3'd2: disp_dat = d[23:20];
        3'd3: disp_dat = d[19:16];
        3'd4: disp_dat = d[15:12];
        3'd5: disp_dat = d[11:8];
        3'd6: disp_dat = d[7:4];
        3'd7: disp_dat = d[3:0];   // самый правый разряд
    endcase

    // В зависимости от count активируем соответствующий разряд
    // Здесь, судя по битам, индикатор с "активным нулём" на разряде:
    // '0' в бите = разряд включён.
    case(count)
        3'd0: dig_r = 8'b0111_1111; // активен разряд 0 (левый)
        3'd1: dig_r = 8'b1011_1111; // активен разряд 1
        3'd2: dig_r = 8'b1101_1111; // активен разряд 2
        3'd3: dig_r = 8'b1110_1111; // активен разряд 3
        3'd4: dig_r = 8'b1111_0111; // активен разряд 4
        3'd5: dig_r = 8'b1111_1011; // активен разряд 5
        3'd6: dig_r = 8'b1111_1101; // активен разряд 6
        3'd7: dig_r = 8'b1111_1110; // активен разряд 7 (правый)
    endcase
end

//--------------------------------------------------------------
// Декодер 4-битного значения в шаблон сегментов
//--------------------------------------------------------------
// seg_r – 8 бит: обычно [dp,g,f,e,d,c,b,a] или подобный порядок.
// Значения 8'hc0, 8'hf9 и т.п. – это "готовые" маски для цифр 0..F.
always @(disp_dat)
begin
    case(disp_dat)
        4'h0: seg_r = 8'hc0;   // отображение '0'
        4'h1: seg_r = 8'hf9;   // '1'
        4'h2: seg_r = 8'ha4;   // '2'
        4'h3: seg_r = 8'hb0;   // '3'
        4'h4: seg_r = 8'h99;   // '4'
        4'h5: seg_r = 8'h92;   // '5'
        4'h6: seg_r = 8'h82;   // '6'
        4'h7: seg_r = 8'hf8;   // '7'
        4'h8: seg_r = 8'h80;   // '8'
        4'h9: seg_r = 8'h90;   // '9'
        4'ha: seg_r = 8'h88;   // 'A'
        4'hb: seg_r = 8'h83;   // 'b'
        4'hc: seg_r = 8'hc6;   // 'C'
        4'hd: seg_r = 8'ha1;   // 'd'
        4'he: seg_r = 8'h86;   // 'E'
        4'hf: seg_r = 8'h8e;   // 'F'
    endcase
end

endmodule
