// Каждый файл Verilog имеет расширение .v (например, filename.v)
// Как и в C/C++, в Verilog также есть однострочные и многострочные комментарии.
// Это однострочный комментарий
/*
   Это многострочный
   комментарий
*/

/*
  Модуль     :   led_water.v
  Создано    : kontakts.ru
  Дата создания : 21-10-2023
  Описание   : Этот модуль моделирует эффект "воды" на LED-ленте с использованием тактового сигнала 50 МГц.
               Светодиоды сдвигаются в каскадном порядке, включаются и выключаются, создавая эффект текущей воды.
*/

module led_water(led, clk); // Модуль является частью аппаратного обеспечения в Verilog. Синтаксис Verilog начинается с "module" и заканчивается "endmodule".

  input clk; // Входной тактовый сигнал, 50 МГц

  output [8:1] led; // Выходной сигнал для 8 LED, представленных 8-битным значением (1 байт)

  reg [8:1] led; // Регистры для хранения состояния LED (8-битное значение)
  reg [24:0] counter; // 25-битный счетчик для управления временем

  // Always блок, срабатывающий на положительном фронте тактового сигнала
  always @(posedge clk) 
  begin
    counter <= counter + 1; // Увеличиваем значение счетчика
    if (counter == 25'd25000000) // Когда счетчик достигает 25 миллионов (для управления временем)
    begin
      led <= led << 1; // Сдвигаем состояние LED влево (эффект каскада)
      counter <= 0; // Сбрасываем счетчик
      if (led == 8'b0000_0000) // Если все LED выключены
        led <= 8'b1111_1111; // Включаем все LED
    end
  end
endmodule

	
