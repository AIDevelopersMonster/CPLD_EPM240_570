// ============================================================
// Имя файла: my_uart_tx.v
// Описание: Модуль передачи данных через UART (RS232). 
//           Обрабатывает передачу данных, синхронизирует их по скорости 
//           передачи и генерирует тактовые сигналы для передачи данных.
//           Модуль управляет состояниями передачи и обработкой байтов данных.
//
// Создано: AIDevelopersMonster
// Репозиторий GitHub: https://github.com/AIDevelopersMonster/CPLD_EPM240_570/
//
// ============================================================

`timescale 1ns / 1ps

module my_uart_tx(
    input clk,            // Входной тактовый сигнал 50MHz
    input rst_n,          // Низкий активный сигнал сброса
    input clk_bps,        // Тактовый сигнал для синхронизации скорости передачи данных
    input [7:0] rx_data, // Принятые 8 бит данных
    input rx_int,         // Сигнал прерывания для начала передачи данных
    output rs232_tx,      // Выходной сигнал передачи данных RS232
    output bps_start      // Сигнал начала передачи данных для синхронизации
);

// Временные регистры для управления прерыванием и состоянием передачи
reg rx_int0, rx_int1, rx_int2;  // Регистры для задержки прерывания
wire neg_rx_int;  // Обнаружение переднего фронта сигнала прерывания

// Сдвиговые регистры для обработки сигнала rx_int
always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        rx_int0 <= 1'b0;
        rx_int1 <= 1'b0;
        rx_int2 <= 1'b0;
    end else begin
        rx_int0 <= rx_int;
        rx_int1 <= rx_int0;
        rx_int2 <= rx_int1;
    end
end

// Обнаружение переднего фронта сигнала rx_int
assign neg_rx_int = ~rx_int1 & rx_int2;  // Когда прерывание изменяется с 0 на 1

//---------------------------------------------------------
// Регистры для хранения данных и управления передачей
reg [7:0] tx_data;  // Данные для передачи
reg bps_start_r;     // Сигнал начала передачи
reg tx_en;           // Включение передачи
reg [3:0] num;       // Счетчик битов для передачи

always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        bps_start_r <= 1'bz;
        tx_en <= 1'b0;
        tx_data <= 8'd0;
    end else if (neg_rx_int) begin  // Начало передачи при получении данных
        bps_start_r <= 1'b1;
        tx_data <= rx_data;  // Передача полученных данных
        tx_en <= 1'b1;       // Включение передачи
    end else if (num == 4'd11) begin  // Завершение передачи (11 бит)
        bps_start_r <= 1'b0;
        tx_en <= 1'b0;
    end
end

assign bps_start = bps_start_r;  // Сигнал начала передачи

//---------------------------------------------------------
// Регистры для передачи данных через RS232
reg rs232_tx_r;  // Регистр для выхода rs232_tx

always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        num <= 4'd0;
        rs232_tx_r <= 1'b1;  // Стартовая линия RS232
    end else if (tx_en) begin  // Если передача активна
        if (clk_bps) begin  // Считывание данных по тактовому сигналу передачи
            num <= num + 1'b1;
            case (num)
                4'd0: rs232_tx_r <= 1'b0;  // Стартовый бит
                4'd1: rs232_tx_r <= tx_data[0];  // Передача бита 0
                4'd2: rs232_tx_r <= tx_data[1];  // Передача бита 1
                4'd3: rs232_tx_r <= tx_data[2];  // Передача бита 2
                4'd4: rs232_tx_r <= tx_data[3];  // Передача бита 3
                4'd5: rs232_tx_r <= tx_data[4];  // Передача бита 4
                4'd6: rs232_tx_r <= tx_data[5];  // Передача бита 5
                4'd7: rs232_tx_r <= tx_data[6];  // Передача бита 6
                4'd8: rs232_tx_r <= tx_data[7];  // Передача бита 7
                4'd9: rs232_tx_r <= 1'b1;  // Стоповый бит
                default: rs232_tx_r <= 1'b1;  // Стоповый бит по умолчанию
            endcase
        end else if (num == 4'd11) num <= 4'd0;  // Сброс счетчика битов
    end
end

assign rs232_tx = rs232_tx_r;  // Выходной сигнал передачи RS232

endmodule
