// Однострочные комментарии в Verilog начинаются с "//".
// Многострочные комментарии начинаются с "/*" и заканчиваются "*/".

/*
  Модуль     : key_led.v
  Автор      : kontakts.ru
  Создан    : 24-10-2023
*/

module key_led( // Модуль с именем 'key_led', который идентифицируется по этому имени. Порты (key, led) передаются в модуль
    input[MSB_reg:LSB_reg]key,   // входной порт 'key', определенный с диапазоном битов от MSB_reg до LSB_reg.
    output[MSB_reg:LSB_reg]led   // выходной порт 'led', определенный с диапазоном битов от MSB_reg до LSB_reg.
);

// Параметры определяют диапазон битов для портов key и led.
parameter MSB_reg = 6;  // Самый старший бит (MSB) для портов key и led
parameter LSB_reg = 1;  // Самый младший бит (LSB) для портов key и led

// Пояснение о соединениях:
// Модули соединяются через порты, которые могут быть входами, выходами или двусторонними (inout).
// Здесь 'key' является входом, а 'led' — выходом.

// Определение регистров:
// 'led_r' хранит состояние светодиодов, и это регистр с шириной 6 бит.
reg[MSB_reg:1]led_r;  // 6-битный регистр для хранения состояния светодиодов
reg[6:LSB_reg]buffer;  // Буферный регистр для временного хранения входного значения 'key'

// Ключевое слово 'assign' используется для присваивания значения выходному порту 'led'.
// Здесь мы присваиваем значение регистра 'led_r' выходному порту 'led'.
assign led = led_r; // Выходной LED присваивается значению, хранящемуся в led_r

// Блок always срабатывает каждый раз, когда значение 'key' изменяется
always @(key) begin
    buffer = key;  // Сохраняем значение 'key' в буфер
    case (buffer)  // Проверяем значение буфера (key)
        6'b111110:               // Если key равно '111110' (key1)
            led_r = 6'b111110;   // Включаем LED1
        6'b111101:               // Если key равно '111101' (key2)
            led_r = 6'b111100;   // Включаем LED1, LED2
        6'b111011:               // Если key равно '111011' (key3)
            led_r = 6'b111000;   // Включаем LED1, LED2, LED3
        6'b110111:               // Если key равно '110111' (key4)
            led_r = 6'b110000;   // Включаем LED1, LED2, LED3, LED4
        6'b101111:               // Если key равно '101111' (key5)
            led_r = 6'b100000;   // Включаем LED1, LED2, LED3, LED4, LED5
        6'b011111:               // Если key равно '011111' (key6)
            led_r = 6'b000000;   // Выключаем все светодиоды (LED1 до LED6)
        default: led_r = 6'b111111; // В случае по умолчанию включаем все светодиоды (LED1 до LED6)
    endcase
end

endmodule  // Конец модуля

/*
Структура модуля Verilog:
1. module <имя_модуля> (
2.   // Определяем все входные и выходные порты
3.   <имя_порта>
4. );
5. 
6.   // Опционально можно объявить параметры
7.   parameter <имя_параметра> = <значение_по_умолчанию>;
8. 
9.   // Завершаем определение портов модуля (входы/выходы)
10.  <направление> <тип_данных> <размер> <имя_порта>;
11. 
12.  // RTL (Register Transfer Level) или структурный код здесь
13. 
14. endmodule

Ключевые концепции Verilog:
1. Ключевые слова такие как module, assign и другие — это зарезервированные слова.
2. Представление бинарных значений в Verilog:
   - 3'b100 означает 3-битное бинарное значение 100.
3. Представление шестнадцатеричных значений в Verilog:
   - 4'h8 означает 8-битное шестнадцатеричное значение 8.
4. Представление октальных значений в Verilog:
   - 4'o10 означает 8-битное октальное значение 10.
5. Представление десятичных значений в Verilog:
   - 4'd8 означает 8-битное десятичное значение 8.

Тип 'Reg' в Verilog используется для определения регистров, которые сохраняют значения и могут удерживать их между тактами.

1. always @(<список_чувствительных_сигналов>) begin  // Блок срабатывает, когда любой из сигналов в списке чувствительности изменяется
2.    // Код, который будет выполнен
3. end
*/
