`timescale 1 ns / 1 ns

/*
  Module     : spidac.v
  Created By : kontakts.ru
  Description: Управление ЦАП TLC5615 по SPI с помощью CPLD EPM240/EPM570.
               Напряжение на выходе ЦАП задаётся положением 4 ползунков ckey[1]..ckey[4].
               Диапазон: от ~0 В до ~5 В (при Vref = 5 В).
*/

module spidac(
    clk,
    Reset,
    dac_sclk,
    DAC_nCS,
    dac_din,
    ckey            // вход — ползунковые переключатели
);
    // -------- ПОРТЫ МОДУЛЯ --------------------------------------
    input            clk;       // Системный тактовый сигнал (например, 50 МГц)
    input            Reset;     // Асинхронный сброс, активный низким уровнем
    output           dac_sclk;  // SPI SCLK для TLC5615
    output           DAC_nCS;   // SPI /CS (chip select), активный низким уровнем
    output           dac_din;   // SPI DIN — последовательные данные для ЦАП
    input  [4:1]     ckey;      // 4 ползунка ckey[1]..ckey[4]

    // ============================================================
    // 1. Делители частоты: получаем более медленный такт для SPI
    //    clk -> clkdiv2 -> clkdiv4 (делим частоту в 4 раза)
    // ============================================================
    reg clkdiv2;
    reg clkdiv4;

    // Делитель на 2
    always @(posedge clk or negedge Reset)
        if (!Reset)
            clkdiv2 <= 1'b0;
        else
            clkdiv2 <= ~clkdiv2;

    // Ещё делитель на 2 (в сумме делим на 4)
    always @(posedge clkdiv2 or negedge Reset)
        if (!Reset)
            clkdiv4 <= 1'b0;
        else
            clkdiv4 <= ~clkdiv4;

    // ============================================================
    // 2. Формирование 10-битного значения для ЦАП из 4 ползунков
    //
    //    ckey[1]..ckey[4] образуют 4-битное число:
    //    level = 0..15  (всего 16 уровней)
    //
    //    Преобразуем:
    //    dac_value = level * 68 ≈ 0..1020  (почти весь 10-битный диапазон)
    //
    //    При Vref = 5 В:
    //      level = 0  → ~0 В
    //      level = 15 → ~4.99 В
    //
    //    Важно: в зависимости от схемотехники ползунков
    //    "ON" может означать 0 или 1. Если направление покажется
    //    "перевёрнутым", можно инвертировать level.
    // ============================================================
    wire [3:0] level = {ckey[4], ckey[3], ckey[2], ckey[1]};  // собираем в правильном порядке

    // Масштабируем 4 бита до 10 бит (0..1020)
    wire [9:0] dac_value = level * 10'd68;

    // ============================================================
    // 3. SPI-логика для TLC5615, 16-битный кадр
    //
    //    TLC5615 ожидает 16 бит:
    //      [15:12] — "don't care" (обычно 0000)
    //      [11:2]  — 10 бит данных D9..D0 (MSB первым)
    //      [1:0]   — "don't care" (обычно 00)
    //
    //    Мы формируем:
    //      shift_reg = {4'b0000, dac_value[9:0], 2'b00}
    // ============================================================
    reg [15:0] shift_reg;   // сдвиговый регистр для SPI-передачи
    reg [4:0]  bit_cnt;     // счётчик бит (0..15)

    // Состояния простой машины состояний
    localparam ST_IDLE = 2'b00;
    localparam ST_LOAD = 2'b01;
    localparam ST_SEND = 2'b10;
    localparam ST_DONE = 2'b11;

    reg [1:0] state;

    // Выходные регистры SPI
    reg sclk_reg;
    reg ncs_reg;

    assign dac_sclk = sclk_reg;       // тактовый сигнал для TLC5615
    assign DAC_nCS  = ncs_reg;        // /CS (active low)
    assign dac_din  = shift_reg[15];  // всегда выдаём старший бит регистра

    // ============================================================
    // 4. Машина состояний SPI:
    //    IDLE -> LOAD -> SEND (16 тактов) -> DONE -> IDLE ...
    // ============================================================
    always @(posedge clkdiv4 or negedge Reset) begin
        if (!Reset) begin
            state     <= ST_IDLE;
            bit_cnt   <= 5'd0;
            shift_reg <= 16'd0;
            sclk_reg  <= 1'b0;
            ncs_reg   <= 1'b1;   // CS неактивен
        end else begin
            case (state)

                //-------------------------------------------------
                // Ожидание — здесь можно вставить паузу или запуск по событию
                //-------------------------------------------------
                ST_IDLE: begin
                    ncs_reg  <= 1'b1;  // отпускаем /CS
                    sclk_reg <= 1'b0;  // линия такта в "0"
                    state    <= ST_LOAD;
                end

                //-------------------------------------------------
                // Загрузка данных в сдвиговый регистр:
                // [15:12] = 0000
                // [11:2]  = dac_value (10 бит)
                // [1:0]   = 00
                //-------------------------------------------------
                ST_LOAD: begin
                    shift_reg <= {4'b0000, dac_value, 2'b00};
                    bit_cnt   <= 5'd0;
                    ncs_reg   <= 1'b0;  // активируем TLC5615 (CS = 0)
                    sclk_reg  <= 1'b0;
                    state     <= ST_SEND;
                end

                //-------------------------------------------------
                // Передача 16 бит по SPI
                //-------------------------------------------------
                ST_SEND: begin
                    // Генерируем тактовый сигнал SCLK
                    sclk_reg <= ~sclk_reg;

                    // Сдвигаем данные и считаем биты на одном из фронтов
                    // Здесь используется "старое" значение sclk_reg:
                    // if (sclk_reg == 1) — значит только что был переход 1->0
                    if (sclk_reg) begin
                        if (bit_cnt == 5'd15) begin
                            state <= ST_DONE; // все 16 бит отправлены
                        end else begin
                            bit_cnt   <= bit_cnt + 1'b1;
                            // Сдвиг влево, на место младшего бита подставляем 0
                            shift_reg <= {shift_reg[14:0], 1'b0};
                        end
                    end
                end

                //-------------------------------------------------
                // Завершение кадра — отпускаем /CS и возвращаемся в IDLE
                //-------------------------------------------------
                ST_DONE: begin
                    ncs_reg  <= 1'b1;   // завершаем передачу
                    sclk_reg <= 1'b0;
                    state    <= ST_IDLE;
                end

                default: begin
                    state <= ST_IDLE;
                end
            endcase
        end
    end

endmodule
