//*******************************************************//
//                Интегральный делитель частоты          //
//*******************************************************//
// Назначение:
//   Делит входную частоту clock во F_DIV раз и формирует
//   выходной сигнал clk_out.
//
//   Параметр F_DIV – коэффициент деления (1..2^n, n = F_DIV_WIDTH).
//   При необходимости изменить частоту на выходе нужно
//   изменить только F_DIV (и при желании F_DIV_WIDTH под его разрядность).
//
//   Если F_DIV чётный – скважность clk_out близка к 50%.
//   Если F_DIV нечётный – используются два счётчика по фронту/спаду,
//   чтобы сделать скважность максимально близкой к 50%.
//
// Пример настроек (если clock = 50 МГц):
//   Нужен 1 кГц  → F_DIV = 50_000
//   Нужен 10 кГц → F_DIV = 5_000
//
// Диаграмма (условно):
//   clock     |--|__|--|__|--|__|--|__|--|__|--|__|
//   clk_p_r   |_____|-----------|_____|-----------| 
//   clk_n_r   ---|_____|-----------|_____|---------
//   clk_out   |________|--------|________|--------|
//
//*******************************************************

module int_div(
    clock,    // входной системный тактовый сигнал
    clk_out   // выходной, разделённый по частоте сигнал
);

// I/O порты
input  clock;     // входной тактовый сигнал
output clk_out;   // выходной сигнал после деления

// Внутренние регистры
reg clk_p_r;                          // делитель по фронту (posedge clock)
reg clk_n_r;                          // делитель по спаду (negedge clock)
reg [F_DIV_WIDTH - 1:0] count_p;      // счётчик для положительного фронта
reg [F_DIV_WIDTH - 1:0] count_n;      // счётчик для отрицательного фронта

// Параметры делителя
parameter F_DIV       = 48000000;     // коэффициент деления <<<<----- менять здесь
parameter F_DIV_WIDTH = 32;           // разрядность счётчиков

// Внутренние флаги
wire full_div_p;      // счётчик по фронту ещё не дошёл до F_DIV - 1
wire half_div_p;      // счётчик по фронту ещё не дошёл до F_DIV/2 - 1
wire full_div_n;      // счётчик по спаду ещё не дошёл до F_DIV - 1
wire half_div_n;      // счётчик по спаду ещё не дошёл до F_DIV/2 - 1

// Условия для сравнения счётчиков
assign full_div_p = (count_p < F_DIV - 1);
assign half_div_p = (count_p < (F_DIV >> 1) - 1);
assign full_div_n = (count_n < F_DIV - 1);
assign half_div_n = (count_n < (F_DIV >> 1) - 1);

// Формирование выходного сигнала
// Если F_DIV = 1 → делитель отключён, clk_out = clock.
// Если F_DIV нечётный → clk_out = clk_p_r & clk_n_r (комбинация двух полупериодов).
// Если F_DIV чётный → используется только clk_p_r.
assign clk_out = (F_DIV == 1) ? 
                 clock : (F_DIV[0] ? (clk_p_r & clk_n_r) : clk_p_r);

//-------------------------------------------------------
// Делитель по положительному фронту clock
//-------------------------------------------------------
always @(posedge clock)
begin
    if (full_div_p)
    begin
        count_p <= count_p + 1'b1;
        if (half_div_p)
            clk_p_r <= 1'b0;          // первая половина периода – низкий уровень
        else
            clk_p_r <= 1'b1;          // вторая половина периода – высокий уровень
    end
    else
    begin
        count_p <= 0;                 // сброс счётчика
        clk_p_r <= 1'b0;
    end
end

//-------------------------------------------------------
// Делитель по отрицательному фронту clock
//-------------------------------------------------------
always @(negedge clock)
begin
    if (full_div_n)
    begin
        count_n <= count_n + 1'b1;
        if (half_div_n)
            clk_n_r <= 1'b0;          // первая половина периода – низкий
        else
            clk_n_r <= 1'b1;          // вторая половина периода – высокий
    end
    else
    begin
        count_n <= 0;                 // сброс счётчика
        clk_n_r <= 1'b0;
    end
end

endmodule
