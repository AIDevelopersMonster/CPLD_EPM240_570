// ------------------------------------------------------------
//  Module     : lcd.v
//  Project    : LCD1602 "HELLO WORLD!" demo для CPLD/FPGA
//  Board      : EPM240 / EPM570 (и подобные, с тактовой частотой ~50 МГц)
//  Created By : kontakts.ru
//  Description: 
//    Простой пример инициализации символьного дисплея LCD1602
//    в 8-битном режиме и вывода строки "HELLO WORLD!" в первую
//    строку дисплея.
//
//    Модуль реализует простой конечный автомат (FSM), который:
//      1) Понижает частоту системного тактового сигнала (делитель).
//      2) Последовательно отправляет команды и данные в контроллер LCD.
//      3) По завершении записи строки оставляет EN в "1", чтобы
//         дисплей оставался инициализированным.
//
//    Репозиторий проекта:
//      https://github.com/AIDevelopersMonster/CPLD_EPM240_570
//
//    Плейлист FPGA / CPLD (YouTube):
//      https://www.youtube.com/playlist?list=PLVoFIRfTAAI7-d_Yk6bNVnj4atUdMxvT5
//
//
// ------------------------------------------------------------


module lcd(clk, rs, rw, en, dat);  

    // clk — входной тактовый сигнал от платы (обычно 50 МГц)
    input clk;  

    // dat — выходные 8-битные данные на LCD1602 (шина D7..D0)
    output [7:0] dat; 

    // rs — выбор регистра LCD:
    //       0 = команда, 1 = данные (символ)
    // rw — режим доступа:
    //       0 = запись в LCD (мы используем только запись)
    // en — строб записи (фронт активирует передачу в LCD)
    output rs, rw, en;
 //tri en; 
  // --------------------------------------------------------
    // Регистры для внутренней логики
    // --------------------------------------------------------
    reg        e;          // Дополнительный бит для формирования сигнала EN
    reg [7:0]  dat;        // Регистр выходных данных на шину D7..D0
    reg        rs;         // Регистр для сигнала RS
    reg [15:0] counter;    // Делитель частоты для получения более медленного такта
    reg [4:0]  current;    // Текущее состояние конечного автомата
    reg [4:0]  next;       // Следующее состояние конечного автомата
    reg        clkr;       // "Замедленный" тактовый сигнал для FSM
    reg [1:0]  cnt;        // Счетчик проходов по инициализации

    // --------------------------------------------------------
    // Коды состояний конечного автомата
    // --------------------------------------------------------
    parameter  set0   = 5'h00; // Команда: начальная настройка (0x30)
    parameter  set1   = 5'h01; // Команда: включение дисплея (0x0C)
    parameter  set2   = 5'h02; // Команда: режим ввода (0x06)
    parameter  set3   = 5'h03; // Команда: очистка дисплея (0x01)

    // Дальше — состояния вывода символов "HELLO WORLD!"
    parameter  dat0   = 5'h04; // 'H'
    parameter  dat1   = 5'h05; // 'E'
    parameter  dat2   = 5'h06; // 'L'
    parameter  dat3   = 5'h07; // 'L'
    parameter  dat4   = 5'h08; // 'O'
    parameter  dat5   = 5'h09; // ' '
    parameter  dat6   = 5'h0A; // 'W'
    parameter  dat7   = 5'h0B; // 'O'
    parameter  dat8   = 5'h0C; // 'R'
    parameter  dat9   = 5'h0D; // 'L'
    parameter  dat10  = 5'h0E; // 'D'
    parameter  dat11  = 5'h10; // '!'
    parameter  nul    = 5'h0F; // Конечное состояние (ожидание)

    // --------------------------------------------------------
    // Делитель частоты: формируем более "медленный" тактовый
    // Для ЖК-дисплея не нужен системный такт 50 МГц, мы его
    // делим, чтобы FSM переключался редко (и выдерживались
    // задержки для LCD).
    // --------------------------------------------------------
    always @(posedge clk) begin
        counter <= counter + 1'b1;

        // Когда счетчик достигает небольшого значения,
        // инвертируем clkr и снова считаем.
        // В реальном проекте значение можно подобрать под
        // реальные тайминги LCD (t > 40 мкс для команд и пр.).
        if (counter == 16'h000F) begin
            clkr    <= ~clkr;
            counter <= 16'h0000;
        end
    end

    // --------------------------------------------------------
    // Конечный автомат управления LCD
    // Срабатывает по "медленному" тактовому сигналу clkr.
    // --------------------------------------------------------
    always @(posedge clkr) begin
        current <= next;   // Переход в следующее состояние

        case (current)
            // ---------------- ИНИЦИАЛИЗАЦИЯ ----------------
            set0: begin
                rs   <= 1'b0;     // Режим команды
                dat  <= 8'h30;    // Функциональная установка (8-битный интерфейс)
                next <= set1;
            end

            set1: begin
                rs   <= 1'b0;
                dat  <= 8'h0C;    // Включить дисплей, курсор выкл., мигание выкл.
                next <= set2;
            end

            set2: begin
                rs   <= 1'b0;
                dat  <= 8'h06;    // Режим ввода: авто-инкремент адреса
                next <= set3;
            end

            set3: begin
                rs   <= 1'b0;
                dat  <= 8'h01;    // Очистка дисплея
                next <= dat0;
            end

            // ---------------- ВЫВОД ТЕКСТА -----------------
            dat0: begin
                rs   <= 1'b1;     // Режим "данные" (символ)
                dat  <= "H";
                next <= dat1;
            end

            dat1: begin
                rs   <= 1'b1;
                dat  <= "E";
                next <= dat2;
            end

            dat2: begin
                rs   <= 1'b1;
                dat  <= "L";
                next <= dat3;
            end

            dat3: begin
                rs   <= 1'b1;
                dat  <= "L";
                next <= dat4;
            end

            dat4: begin
                rs   <= 1'b1;
                dat  <= "O";
                next <= dat5;
            end

            dat5: begin
                rs   <= 1'b1;
                dat  <= " ";
                next <= dat6;
            end

            dat6: begin
                rs   <= 1'b1;
                dat  <= "W";
                next <= dat7;
            end

            dat7: begin
                rs   <= 1'b1;
                dat  <= "O";
                next <= dat8;
            end

            dat8: begin
                rs   <= 1'b1;
                dat  <= "R";
                next <= dat9;
            end

            dat9: begin
                rs   <= 1'b1;
                dat  <= "L";
                next <= dat10;
            end

            dat10: begin
                rs   <= 1'b1;
                dat  <= "D";
                next <= dat11;
            end

            dat11: begin
                rs   <= 1'b1;
                dat  <= "!";
                next <= nul;
            end

            // ---------------- ФИНАЛЬНОЕ СОСТОЯНИЕ -----------
            nul: begin
                rs  <= 1'b0;
                dat <= 8'h00;   // Можно отправлять "пустую" команду

                // cnt — счетчик повторов инициализации.
                // Пока меньше 2 — снова запускаем инициализацию.
                // Потом останавливаемся в текущем состоянии.
                if (cnt != 2'h2) begin
                    e    <= 1'b0;
                    next <= set0;   // Повторить инициализацию
                    cnt  <= cnt + 1'b1;
                end
                else begin
                    next <= nul;    // Остаемся здесь
                    e    <= 1'b1;   // Защелкиваем EN
                end
            end

            // На всякий случай — возврат к началу
            default: begin
                next <= set0;
            end
        endcase
    end

    // --------------------------------------------------------
    // Формирование выходных сигналов
    // --------------------------------------------------------
    assign en = clkr | e;  // EN активен при тактовой активности или в финале
    assign rw = 1'b0;      // Всегда пишем в дисплей

endmodule