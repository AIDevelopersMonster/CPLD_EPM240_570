// Одиночный комментарий в Verilog начинается с // 
// Многострочные комментарии начинаются с /* и заканчиваются на */

//------------------------------------------------------------------
// Модуль: sled.v
// Описание: Модуль для управления 7-сегментным дисплеем. Используется 
// для отображения чисел от 0 до 15 (в формате 4-битного числа) на дисплее.
// Создано: kontakts.ru
// Дата создания: 26-10-2023
//------------------------------------------------------------------

module sled(seg, dig, clock); // Объявление модуля с портами

    input clock;               // Вход: тактовый сигнал (clock)
    output [7:0] seg;          // Выход: 8 бит для управления сегментами дисплея
    output [7:0] dig;          // Выход: 8 бит для управления цифрами дисплея

    reg [7:0] seg;             // Регистр для хранения текущего состояния сегментов
    reg [7:0] dig;             // Регистр для хранения текущего состояния разрядов
    reg [3:0] disp_dat;        // Регистр для хранения данных, которые отображаются на дисплее
    reg [36:0] count;          // Регистр для счётчика, чтобы создавать задержки

    // Основной блок, который увеличивает счётчик на каждом фронте тактового сигнала
    always @ (posedge clock) begin
        count = count + 1'b1;    // Увеличиваем счётчик на 1
        dig = 8'b00000000;        // Очистка дисплея (по умолчанию все разряды выключены)
    end

    // Этот блок срабатывает по изменению 24-го бита счётчика
    always @ (count[24]) begin
        // Используется 4 старших бита для отображения чисел от 0 до 15
        disp_dat = {count[28:25]}; // disp_dat будет содержать значения от 0000 до 1111 (от 0 до 15)
    end

    // Блок, который управляет отображением числа на дисплее в зависимости от disp_dat
    always @ (disp_dat) begin
        // В зависимости от значения disp_dat выбираем, какие сегменты включить для отображения числа
        case (disp_dat)
            4'h0 : seg = 8'hc0; // "0"
            4'h1 : seg = 8'hf9; // "1"
            4'h2 : seg = 8'hA4; // "2"
            4'h3 : seg = 8'hb0; // "3"
            4'h4 : seg = 8'h99; // "4"
            4'h5 : seg = 8'h92; // "5"
            4'h6 : seg = 8'h82; // "6"
            4'h7 : seg = 8'hf8; // "7"
            4'h8 : seg = 8'h80; // "8"
            4'h9 : seg = 8'h90; // "9"
            4'ha : seg = 8'h88; // "a"
            4'hb : seg = 8'h83; // "b"
            4'hc : seg = 8'hc6; // "c"
            4'hd : seg = 8'ha1; // "d"
            4'he : seg = 8'h86; // "e"
            4'hf : seg = 8'h8e; // "f"
        endcase
    end

endmodule

