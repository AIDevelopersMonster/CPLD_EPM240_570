`timescale 1ns / 1ps

module speed_select(
				clk,rst_n,
				bps_start,clk_bps
			);

input clk;	        // Тактовый сигнал 50 МГц
input rst_n;	    // Сброс, активный низкий уровень
input bps_start;	// Старт работы делителя: 1 — идёт передача, нужно формировать clk_bps
output clk_bps;	    // Тактовый импульс для UART: высокий уровень в момент выборки следующего бита

/*
parameter 		bps9600 	= 5207,	// делитель для скорости 9600 bps
			 	bps19200 	= 2603,	// делитель для скорости 19200 bps
				bps38400 	= 1301,	// делитель для скорости 38400 bps
				bps57600 	= 867,	// делитель для скорости 57600 bps
				bps115200	= 433;	// делитель для скорости 115200 bps

parameter 		bps9600_2 	= 2603,
				bps19200_2	= 1301,
				bps38400_2	= 650,
				bps57600_2	= 433,
				bps115200_2 = 216;  
*/

	// Ниже выбраны конкретные значения делителей под нужную скорость UART.
	// При желании скорость можно изменить, пересчитав BPS_PARA и BPS_PARA_2.
`define		BPS_PARA		5207	// Делитель для скорости 9600 bps (полный период)
`define 	BPS_PARA_2		2603	// Половина периода для 9600 bps — момент выборки бита

reg[12:0] cnt;			// Делитель частоты (счётчик для формирования clk_bps)
reg clk_bps_r;			// Регистр формирования тактового импульса clk_bps

//----------------------------------------------------------
reg[2:0] uart_ctrl;	// Зарезервирован под выбор режима UART (сейчас не используется)
//----------------------------------------------------------

always @ (posedge clk or negedge rst_n)
	if(!rst_n) cnt <= 13'd0;
	else if((cnt == `BPS_PARA) || !bps_start) cnt <= 13'd0;	// При достижении максимума или при остановке bps_start — сброс счётчика
	else cnt <= cnt+1'b1;			// В остальных случаях счётчик просто увеличивается

always @ (posedge clk or negedge rst_n)
	if(!rst_n) clk_bps_r <= 1'b0;
	else if(cnt == `BPS_PARA_2) clk_bps_r <= 1'b1;	// clk_bps_r в 1 только в середине периода — момент выборки бита данных
	else clk_bps_r <= 1'b0;

assign clk_bps = clk_bps_r;

endmodule
