// ============================================================
// Имя файла: speed_select.v
// Описание: Модуль для генерации тактового сигнала с заданной скоростью
//           (baud rate). Модуль принимает сигнал начала передачи данных
//           и генерирует тактовый сигнал для синхронизации передачи данных.
//           Поддерживает различные скорости передачи данных.
//
// Создано: AIDevelopersMonster
// Репозиторий GitHub: https://github.com/AIDevelopersMonster/CPLD_EPM240_570/
//
// ============================================================

`timescale 1ns / 1ps

module speed_select(
    input clk,        // Входной тактовый сигнал 50MHz
    input rst_n,      // Низкий активный сигнал сброса
    input bps_start,  // Сигнал начала передачи данных
    output clk_bps    // Выходной тактовый сигнал для передачи данных
);

// Параметры для различных скоростей передачи данных (baud rates)
`define BPS_PARA     5207    // Для скорости 9600bps
`define BPS_PARA_2   2603    // Для скорости 9600bps (вторая часть для делителя)

reg [12:0] cnt;        // Счётчик для отслеживания тактов
reg clk_bps_r;         // Внутренний тактовый сигнал для передачи данных

//----------------------------------------------------------
// Регистры для управления состоянием UART
//----------------------------------------------------------

always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        cnt <= 13'd0;  // Сброс счётчика при сбросе
    end else if ((cnt == `BPS_PARA) || !bps_start) begin
        cnt <= 13'd0;  // Если счётчик достигает заданного значения, сбрасываем
    end else begin
        cnt <= cnt + 1'b1;  // Увеличиваем счётчик при каждом такте
    end
end

always @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        clk_bps_r <= 1'b0;  // Сброс тактового сигнала при сбросе
    end else if (cnt == `BPS_PARA_2 && bps_start) begin
        clk_bps_r <= 1'b1;  // Генерация тактового сигнала для передачи данных
    end else begin
        clk_bps_r <= 1'b0;  // Отключение тактового сигнала, если счётчик не равен нужному значению
    end
end

assign clk_bps = clk_bps_r;  // Выходной тактовый сигнал

endmodule
