//--------------------------------------------------------------------------------------------------
// step_moto.v — управление шаговым двигателем (8-состояний, полушаговый режим)
//
// Функции модуля:
// - Делитель частоты от системного тактового сигнала clk.
// - Формирование последовательности сигналов StepDrive[3:0] для управления 4 обмотками двигателя.
// - Направление вращения задаётся сигналом Dir.
// - Пуск/останов вращения — сигналом StepEnable.
// - Асинхронный сброс rst (активный низкий уровень).
//
// Пример: при StepLockOut = 200000 и частоте clk ≈ 50 МГц
//         частота шагов ≈ 50e6 / 200000 ≈ 250 Гц.
//--------------------------------------------------------------------------------------------------

module step_moto (
    StepDrive,   // 4 выхода на ключи / драйверы обмоток шагового двигателя
    clk,         // системный тактовый сигнал (например, 50 МГц)
    Dir,         // направление вращения: 1 — вперёд, 0 — назад
    StepEnable,  // разрешение вращения: 1 — запуск, 0 — останов
    rst          // асинхронный сброс (активный низкий уровень)
);

    input clk;
    input Dir;
    input StepEnable;
    input rst;

    output [3:0] StepDrive;
    reg    [3:0] StepDrive;   // текущий шаблон управления обмотками

    reg [2:0]  state;         // номер текущего шага (0..7)
    reg [31:0] StepCounter = 32'b0;  // счётчик для деления частоты
    // Параметр делителя частоты — задаёт скорость вращения двигателя
    parameter [31:0] StepLockOut = 32'd200000; // ≈250 Гц при 50 МГц
    reg InternalStepEnable;   // внутренний флаг, фиксирующий запуск

    // Асинхронный сброс по низкому уровню rst и логика счётчика/состояний
    always @(posedge clk or negedge rst)
    begin
        // rst = 0 -> сбрасываем все регистры
        if (!rst) begin
            StepDrive          <= 4'b0000;
            state              <= 3'b000;
            StepCounter        <= 32'b0;
            InternalStepEnable <= 1'b0;
        end
        else begin
            // Если пришла команда на старт — запоминаем её
            if (StepEnable == 1'b1)
                InternalStepEnable <= 1'b1;

            // Делитель частоты: считаем до StepLockOut
            StepCounter <= StepCounter + 32'b1;
            if (StepCounter >= StepLockOut) begin
                StepCounter <= 32'b0;

                // Если внутренний флаг разрешён — делаем шаг
                if (InternalStepEnable == 1'b1) begin
                    // Обновляем внутренний флаг по текущему входу StepEnable
                    // (при StepEnable = 0 двигатель остановится после текущего шага)
                    InternalStepEnable <= StepEnable;

                    // Выбор направления: вперёд / назад
                    if (Dir == 1'b1)
                        state <= state + 3'b001;   // шаг вперёд
                    else
                        state <= state - 3'b001;   // шаг назад

                    // Таблица состояний для управления обмотками
                    // Последовательность даёт полушаговый режим (8 состояний)
                   case (state)
                        3'b000: StepDrive <= 4'b0001; // Обмотка 1
                        3'b001: StepDrive <= 4'b0011; // 1 + 2
                        3'b010: StepDrive <= 4'b0010; // Обмотка 2
                        3'b011: StepDrive <= 4'b0110; // 2 + 3
                        3'b100: StepDrive <= 4'b0100; // Обмотка 3
                        3'b101: StepDrive <= 4'b1100; // 3 + 4
                        3'b110: StepDrive <= 4'b1000; // Обмотка 4
                        3'b111: StepDrive <= 4'b1001; // 4 + 1
                        default: StepDrive <= 4'b0000;
                    endcase



                end
            end
        end
    end

endmodule
